// Copyright (2019-2022) Paul Scherrer Institute
// SPDX-License-Identifier: CERN-OHL-S-2.0

`timescale 1 ps / 1 ps

module action_wrapper
   (  input           ap_clk,
      input           ap_rst_n,
      input           refclk300_n,
      input           refclk300_p,
      input           gt_ref_clk_n,
      input           gt_ref_clk_p,
      input           gt_rx_gt_port_0_n,
      input           gt_rx_gt_port_0_p,
      input           gt_rx_gt_port_1_n,
      input           gt_rx_gt_port_1_p,
      input           gt_rx_gt_port_2_n,
      input           gt_rx_gt_port_2_p,
      input           gt_rx_gt_port_3_n,
      input           gt_rx_gt_port_3_p,
      output          gt_tx_gt_port_0_n,
      output          gt_tx_gt_port_0_p,
      output          gt_tx_gt_port_1_n,
      output          gt_tx_gt_port_1_p,
      output          gt_tx_gt_port_2_n,
      output          gt_tx_gt_port_2_p,
      output          gt_tx_gt_port_3_n,
      output          gt_tx_gt_port_3_p,
      output          interrupt,
      input           interrupt_ack,
      output [8:0]    interrupt_ctx,
      output [63:0]   interrupt_src,
      output          user_led_a0,
      output          user_led_a1,
      output          user_led_g0,
      output          user_led_g1,

      input           uc_avr_rx,
      output          uc_avr_tx,
      input           uc_avr_ck,

      inout           qsfpdd_scl,
      inout           qsfpdd_sda,
      input           qsfpdd_modprs,
      output [63:0]   m_axi_host_mem_araddr,
      output [1:0]    m_axi_host_mem_arburst,
      output [3:0]    m_axi_host_mem_arcache,
      output [3:0]    m_axi_host_mem_arid,
      output [7:0]    m_axi_host_mem_arlen,
      output [0:0]    m_axi_host_mem_arlock,
      output [2:0]    m_axi_host_mem_arprot,
      output [3:0]    m_axi_host_mem_arqos,
      input           m_axi_host_mem_arready,
      output [3:0]    m_axi_host_mem_arregion,
      output [2:0]    m_axi_host_mem_arsize,
      output [8:0]    m_axi_host_mem_aruser,
      output          m_axi_host_mem_arvalid,
      output [63:0]   m_axi_host_mem_awaddr,
      output [1:0]    m_axi_host_mem_awburst,
      output [3:0]    m_axi_host_mem_awcache,
      output [3:0]    m_axi_host_mem_awid,
      output [7:0]    m_axi_host_mem_awlen,
      output [0:0]    m_axi_host_mem_awlock,
      output [2:0]    m_axi_host_mem_awprot,
      output [3:0]    m_axi_host_mem_awqos,
      input           m_axi_host_mem_awready,
      output [3:0]    m_axi_host_mem_awregion,
      output [2:0]    m_axi_host_mem_awsize,
      output [8:0]    m_axi_host_mem_awuser,
      output          m_axi_host_mem_awvalid,
      input [3:0]     m_axi_host_mem_bid,
      output          m_axi_host_mem_bready,
      input [1:0]     m_axi_host_mem_bresp,
      input [8:0]     m_axi_host_mem_buser,
      input           m_axi_host_mem_bvalid,
      input [1023:0]  m_axi_host_mem_rdata,
      input [3:0]     m_axi_host_mem_rid,
      input           m_axi_host_mem_rlast,
      output          m_axi_host_mem_rready,
      input [1:0]     m_axi_host_mem_rresp,
      input [8:0]     m_axi_host_mem_ruser,
      input           m_axi_host_mem_rvalid,
      output [1023:0] m_axi_host_mem_wdata,
      output          m_axi_host_mem_wlast,
      input           m_axi_host_mem_wready,
      output [127:0]  m_axi_host_mem_wstrb,
      output [8:0]    m_axi_host_mem_wuser,
      output          m_axi_host_mem_wvalid,

      input [31:0]    s_axi_ctrl_reg_araddr,
      input [2:0]     s_axi_ctrl_reg_arprot,
      output          s_axi_ctrl_reg_arready,
      input           s_axi_ctrl_reg_arvalid,
      input [31:0]    s_axi_ctrl_reg_awaddr,
      input [2:0]     s_axi_ctrl_reg_awprot,
      output          s_axi_ctrl_reg_awready,
      input           s_axi_ctrl_reg_awvalid,
      input           s_axi_ctrl_reg_bready,
      output [1:0]    s_axi_ctrl_reg_bresp,
      output          s_axi_ctrl_reg_bvalid,
      output [31:0]   s_axi_ctrl_reg_rdata,
      input           s_axi_ctrl_reg_rready,
      output [1:0]    s_axi_ctrl_reg_rresp,
      output          s_axi_ctrl_reg_rvalid,
      input [31:0]    s_axi_ctrl_reg_wdata,
      output          s_axi_ctrl_reg_wready,
      input [3:0]     s_axi_ctrl_reg_wstrb,
      input           s_axi_ctrl_reg_wvalid
      );

  assign m_axi_host_mem_awuser = 0;
  assign m_axi_host_mem_aruser = 0;
  assign m_axi_host_mem_arlock = 0;
  assign m_axi_host_mem_awlock = 0;
  assign m_axi_host_mem_arregion = 0;
  assign m_axi_host_mem_awregion = 0;
  assign m_axi_host_mem_arqos = 0;
  assign m_axi_host_mem_awqos = 0;
  assign interrupt = 0;
  assign interrupt_src = 0;
  assign interrupt_ctx = 0;

  wire qsfpdd_scl_i;
  wire qsfpdd_scl_o;
  wire qsfpdd_scl_t;
  wire qsfpdd_sda_i;
  wire qsfpdd_sda_o;
  wire qsfpdd_sda_t;

  action action_i
       (.ap_clk(ap_clk),
        .ap_rst_n(ap_rst_n),
        .ref300_clk_n                ( refclk300_n                   ),
        .ref300_clk_p                ( refclk300_p                   ),
        .gt_ref_clk_n                ( gt_ref_clk_n                  ),
        .gt_ref_clk_p                ( gt_ref_clk_p                  ),
        .gt_100g_grx_n               ({gt_rx_gt_port_3_n,gt_rx_gt_port_2_n,gt_rx_gt_port_1_n,gt_rx_gt_port_0_n}),
        .gt_100g_grx_p               ({gt_rx_gt_port_3_p,gt_rx_gt_port_2_p,gt_rx_gt_port_1_p,gt_rx_gt_port_0_p}),
        .gt_100g_gtx_n               ({gt_tx_gt_port_3_n,gt_tx_gt_port_2_n,gt_tx_gt_port_1_n,gt_tx_gt_port_0_n}),
        .gt_100g_gtx_p               ({gt_tx_gt_port_3_p,gt_tx_gt_port_2_p,gt_tx_gt_port_1_p,gt_tx_gt_port_0_p}),
        .qsfpdd_modprs               ( qsfpdd_modprs                 ),

        .m_axi_host_mem_araddr       ( m_axi_host_mem_araddr),
        .m_axi_host_mem_arburst      ( m_axi_host_mem_arburst),
        .m_axi_host_mem_arcache      ( m_axi_host_mem_arcache),
        .m_axi_host_mem_arid         ( m_axi_host_mem_arid),
        .m_axi_host_mem_arlen        ( m_axi_host_mem_arlen),
        .m_axi_host_mem_arprot       ( m_axi_host_mem_arprot),
        .m_axi_host_mem_arready      ( m_axi_host_mem_arready),
        .m_axi_host_mem_arsize       ( m_axi_host_mem_arsize),
        .m_axi_host_mem_arvalid      ( m_axi_host_mem_arvalid),
        .m_axi_host_mem_awaddr       ( m_axi_host_mem_awaddr),
        .m_axi_host_mem_awburst      ( m_axi_host_mem_awburst),
        .m_axi_host_mem_awcache      ( m_axi_host_mem_awcache),
        .m_axi_host_mem_awid         ( m_axi_host_mem_awid),
        .m_axi_host_mem_awlen        ( m_axi_host_mem_awlen),
        .m_axi_host_mem_awprot       ( m_axi_host_mem_awprot),
        .m_axi_host_mem_awready      ( m_axi_host_mem_awready),
        .m_axi_host_mem_awsize       ( m_axi_host_mem_awsize),
        .m_axi_host_mem_awvalid      ( m_axi_host_mem_awvalid),
        .m_axi_host_mem_bready       ( m_axi_host_mem_bready),
        .m_axi_host_mem_bresp        ( m_axi_host_mem_bresp),
        .m_axi_host_mem_bvalid       ( m_axi_host_mem_bvalid),
        .m_axi_host_mem_rdata        ( m_axi_host_mem_rdata),
        .m_axi_host_mem_rlast        ( m_axi_host_mem_rlast),
        .m_axi_host_mem_rready       ( m_axi_host_mem_rready),
        .m_axi_host_mem_rresp        ( m_axi_host_mem_rresp),
        .m_axi_host_mem_rvalid       ( m_axi_host_mem_rvalid),
        .m_axi_host_mem_wdata        ( m_axi_host_mem_wdata),
        .m_axi_host_mem_wlast        ( m_axi_host_mem_wlast),
        .m_axi_host_mem_wready       ( m_axi_host_mem_wready),
        .m_axi_host_mem_wstrb        ( m_axi_host_mem_wstrb),
        .m_axi_host_mem_wvalid       ( m_axi_host_mem_wvalid),
        .s_axi_ctrl_reg_araddr       ( s_axi_ctrl_reg_araddr),
        .s_axi_ctrl_reg_arprot       ( s_axi_ctrl_reg_arprot),
        .s_axi_ctrl_reg_arready      ( s_axi_ctrl_reg_arready),
        .s_axi_ctrl_reg_arvalid      ( s_axi_ctrl_reg_arvalid),
        .s_axi_ctrl_reg_awaddr       ( s_axi_ctrl_reg_awaddr),
        .s_axi_ctrl_reg_awprot       ( s_axi_ctrl_reg_awprot),
        .s_axi_ctrl_reg_awready      ( s_axi_ctrl_reg_awready),
        .s_axi_ctrl_reg_awvalid      ( s_axi_ctrl_reg_awvalid),
        .s_axi_ctrl_reg_bready       ( s_axi_ctrl_reg_bready),
        .s_axi_ctrl_reg_bresp        ( s_axi_ctrl_reg_bresp),
        .s_axi_ctrl_reg_bvalid       ( s_axi_ctrl_reg_bvalid),
        .s_axi_ctrl_reg_rdata        ( s_axi_ctrl_reg_rdata),
        .s_axi_ctrl_reg_rready       ( s_axi_ctrl_reg_rready),
        .s_axi_ctrl_reg_rresp        ( s_axi_ctrl_reg_rresp),
        .s_axi_ctrl_reg_rvalid       ( s_axi_ctrl_reg_rvalid),
        .s_axi_ctrl_reg_wdata        ( s_axi_ctrl_reg_wdata),
        .s_axi_ctrl_reg_wready       ( s_axi_ctrl_reg_wready),
        .s_axi_ctrl_reg_wstrb        ( s_axi_ctrl_reg_wstrb),
        .s_axi_ctrl_reg_wvalid       ( s_axi_ctrl_reg_wvalid),

        .uc_avr_rx                   ( uc_avr_rx),
        .uc_avr_tx                   ( uc_avr_tx),
        .uc_avr_ck                   ( uc_avr_ck),

        .user_led_a0                 ( user_led_a0),
        .user_led_a1                 ( user_led_a1),
        .user_led_g0                 ( user_led_g0),
        .user_led_g1                 ( user_led_g1));

endmodule
